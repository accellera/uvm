//Common testbench for these test case
//3.4        Advanced phase control 5
//  3.4.1         Killing phases. 5
//  3.4.2         Rerunning phases. 5
//  3.4.3         Fast-forwarding. 5

`include "top_uvc.svh"
`include "bot_uvc.svh"
`include "my_seqr.svh"

`include "test_base.svh"