package mem_agent;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "mem_seq_item.svh"
  `include "mem_agent.svh"

endpackage
