// $Id: uvm_tlm.svh,v 1.13 2009/05/01 14:34:38 redelman Exp $
//----------------------------------------------------------------------
//   Copyright 2007-2009 Mentor Graphics Corporation
//   Copyright 2007-2009 Cadence Design Systems, Inc.
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------

`include "uvm_tlm/uvm_tlm_ifs.svh"
`include "uvm_tlm/sqr_ifs.svh"
`include "base/uvm_port_base.svh"

`include "uvm_tlm/uvm_tlm_imps.svh"

`include "uvm_tlm/uvm_imps.svh"
`include "uvm_tlm/uvm_ports.svh"
`include "uvm_tlm/uvm_exports.svh"

`include "uvm_tlm/uvm_tlm_fifo_base.svh"
`include "uvm_tlm/uvm_tlm_fifos.svh"
`include "uvm_tlm/uvm_tlm_req_rsp.svh"

`include "uvm_tlm/sqr_connections.svh"

