module dummy;
endmodule
