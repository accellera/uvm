// $Id: //dvt/vtech/dev/main/avm/cookbook/09_modules/tb_sv/tb_transactor_pkg.sv#2 $
//----------------------------------------------------------------------
//   Copyright 2005-2007 Mentor Graphics Corporation
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------

package hfpb_pkg;

  import uvm_pkg::*;

  `include "hfpb_vif.svh" 
  `include "hfpb_transaction.svh"  
  `include "hfpb_seq_items.svh"  
  `include "hfpb_mapper.svh"
  `include "hfpb_driver.svh"
  `include "hfpb_master.svh"
  `include "hfpb_slave.svh"
  `include "hfpb_responder.svh"
  `include "hfpb_monitor.svh"
  `include "hfpb_coverage.svh"
  `include "hfpb_talker.svh"
  `include "hfpb_sequencer.svh"
  `include "hfpb_agent.svh"
  
endpackage
