//------------------------------------------------------------------------------
// Copyright 2008 Mentor Graphics Corporation
// All Rights Reserved Worldwide
// 
// Licensed under the Apache License, Version 2.0 (the "License"); you may
// not use this file except in compliance with the License.  You may obtain
// a copy of the License at
// 
//        http://www.apache.org/licenses/LICENSE-2.0
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS, WITHOUT
// WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.  See the
// License for the specific language governing permissions and limitations
// under the License.
//------------------------------------------------------------------------------

`ifndef UVM_VMM_PKG_SV
`define UVM_VMM_PKG_SV

`define VMM_UVM_INTEROP
`define VMM_IN_PACKAGE

`include "uvm_pkg.sv"
import uvm_pkg::*;
`include "vmm.sv"

`include "avt_adapters.sv"
import avt_interop_pkg::*;

`endif // UVM_VMM_PKG_SV
