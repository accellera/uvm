//
//----------------------------------------------------------------------
//   Copyright 2013 Freescale Semiconductor, Inc.
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------

`ifndef UVM_ITEM_ALLOCATOR__SVH
`define UVM_ITEM_ALLOCATOR__SVH


//------------------------------------------------------------------------------
//
// CLASS: uvm_converter #(T,I)
//
//------------------------------------------------------------------------------
// A base class for conversion between object representation and integral
// representation.
// This class is virtual and its virtual functions are not implemented.
// They need to be implemented by derived classes.
//------------------------------------------------------------------------------
virtual class uvm_converter#(type T = int, type I = int);
  // Function: serialize
  //
  // Returns integral representation for the given object representation
  virtual  function I serialize(T object);
  endfunction: serialize

  // Function: deserialize
  //
  // Returns object representation for the given integral representation
  virtual function T deserialize(I item);
  endfunction: deserialize
endclass: uvm_converter

//------------------------------------------------------------------------------
//
// CLASS: uvm_simple_converter #(I)
//
//------------------------------------------------------------------------------
// A simple implementation of uvm_converter when object representation is
// equal to integral representation.
//------------------------------------------------------------------------------
class uvm_simple_converter#(type I = int) extends uvm_converter#(I,I);
  // Function: serialize
  //
  // Returns integral representation for the given object representation
  virtual function I serialize(I object);
    return object;
  endfunction: serialize

  // Function: deserialize
  //
  // Returns object representation for the given integral representation
  virtual function I deserialize(I item);
    return item;
  endfunction: deserialize
endclass: uvm_simple_converter


//------------------------------------------------------------------------------
//
// CLASS: uvm_item_alloc_policy #(T,I)
//
//------------------------------------------------------------------------------
// A base class for allocation policy.
//
// An instance of this class is randomized to obtain an allocated item.
// Constraint which does not allow to allocate taken items it provided
// in this class.
//
// This class can be extended to provide additional constraints
// on the allocated item, as validy constraint, since the range of valid items
// is unknown in the generic base class.
//------------------------------------------------------------------------------

class uvm_item_alloc_policy #(type T=longint unsigned, type I=longint unsigned);
  // Parameter: T
  //
  // Specifies the type for object representation of allocated item.
  //

  // Parameter: I
  //
  // Specifies the integral type used for randomization
  //

  uvm_converter#(T,I) converter;

  function new();  
  endfunction: new

  // Variable: item
  //
  // ~item~ is the random member of this class
  // random allocation is done by providing a value to this member.
  // 
  rand I item;

  
  // Variable: object
  //
  // Object representation of allocated item
  // Set in post_randomize();
  //
  T object;
  
  // Variable: in_use
  //
  // Stores all items previously allocated and not released
  // (integral representation)
  //
  I in_use[$];

  // Constraint: not_taken
  //
  // Ensures that sure previously allocated items cannot be selected
  // in the new allocation
  constraint not_taken
  {
    foreach (in_use[i])
    item != in_use[i];
  }

  // A validity constraint (if needed) should be added in any derived
  // classes, as we do not know the list/range of valid items


  // Function: post_randomize
  //
  // Sets the object representation of the allocated object
  function void post_randomize();
    if (converter == null) begin
      `uvm_error("ITEM_ALLOCATOR", "coverter is not set. can not randomize the object")
      return;
    end
    
    object = converter.deserialize(item);
  endfunction: post_randomize
     
endclass: uvm_item_alloc_policy


//------------------------------------------------------------------------------
// Class: uvm_item_allocator
//------------------------------------------------------------------------------
// Main allocator for specific item type
//------------------------------------------------------------------------------
class uvm_item_allocator #(type T=longint unsigned, type I=longint unsigned);

  uvm_item_alloc_policy#(T, I) alloc_policy;

  string  key;  // Used to access global (C side) DB; 
  // If key is empty, global DB is not used and allocator works in local mode

  // Variable: is_local
  //
  // is_local == 0 means that the allocation data base is stored on Verilog side
  // is_local == 1 means that the allocation data base is stored on C side
  bit     is_local;

  // Function: new
  //
  // Creates a new allocator object with the given  ~name~.
  // ~key~ is used to access external allocation database.
  // If ~key~ is empty, the allocation database is stored locally
  // on Verilog side.
  function new(string name, string key = "" );
    this.key = key;
    this.is_local = (key == "");
  endfunction: new
  
  // Variable: in_use
  //
  // Stores all items previously allocated and not released
  // (integral representation)
  //
  protected I in_use[$];


  // Task API

  // Task: lock
  //
  // Locks the external database.
  // Waits if the database is currently locked.
  task lock();
    svdpi_lock_taken_list(key);
  endtask: lock
 
  // Function: unlock
  //
  // removed lock from the external database
  function void unlock();
    svdpi_unlock_taken_list(key);
  endfunction: unlock
  

  // Task: reserve_item_t
  //
  // Reserve specified item -- ~item_to_reserve~.
  //
  // output ~result~ is set to 1 if the item was successfully reserved
  // and to 0 otherwise.

  task reserve_item_t(T item_to_reserve, output bit result);
    lock();
    result = reserve_item(item_to_reserve, 1);
    unlock();
  endtask: reserve_item_t


  // Task: request_item_t
  //
  // Request and reserve an ~item~ according to the specified ~alloc~ policy
  //
  // Output ~result~ is set to 1 if the item was successfully reserved
  // and 0 if otherwise.
  // output ~item~ is set to the allocated item, if allocation was successfull

  task request_item_t(uvm_item_alloc_policy#(T, I) alloc, 
                    output T item, output bit result);
    lock();
    result = request_item(alloc,item,1);
    unlock();
  endtask: request_item_t
 
  // Task: release_item_t
  //
  // Release specified ~object~.
  //
  task release_item_t(T object);
    lock();
    release_item(object,1);
    unlock();
  endtask: release_item_t
  
  // Task: release_all_items_t
  //
  // Release all currenly allocated items
  //
  task release_all_items_t();
    lock();
    release_all_items(1);
    unlock();
  endtask: release_all_items_t


  // Function API


  protected function void import_in_use(bit external_lock = 0);
    // check that size of I is <= 64 bits
    if (!is_local) begin
      int unsigned size;
      longint db[];
      if (!external_lock) begin
        if (svdpi_try_lock_taken_list(key) != 0) // Unsuccessful lock
          `uvm_fatal("ITEM_ALLOCATOR", "lock is not available and function version is called")
      end
      size = svdpi_get_num_taken(key);
      if (size > 0) begin
        db = new[size];
        svdpi_get_taken_list(key,size,db);
        in_use = {};

        for (int unsigned index = 0; index != size; ++index)
        begin
          I value;
          value = db[index];
          in_use.push_back(value);
        end
      end
      else
        in_use = {};
    end
  endfunction: import_in_use

  protected function void export_in_use(bit external_lock = 0); 
    // check that size of I is <= 64 bits
    if (!is_local) begin
      longint db[];
      if (in_use.size() > 0) begin
        db = new[in_use.size()];
        for (int unsigned index = 0; index != in_use.size(); ++index)
          db[index] = in_use[index];
      end
      svdpi_set_taken_list(key,in_use.size(),db);
      if (!external_lock)
        svdpi_unlock_taken_list(key);
    end
  endfunction: export_in_use
  

  protected function void done_in_use(bit external_lock = 0);
    if (!is_local && !external_lock)
       svdpi_unlock_taken_list(key);
  endfunction: done_in_use

  protected function void start_in_use(bit external_lock = 0);
    if (!is_local && !external_lock)
       begin
         if (svdpi_try_lock_taken_list(key) != 0) // Unsuccessful lock
          `uvm_fatal("ITEM_ALLOCATOR", "Lock is not available and function version of DB access has been called.  Cannot wait for lock")
       end
  endfunction: start_in_use


  // Function: can_reserve
  //
  // Check if the specified ~item_to_reserve~ can be reserved.
  // Returns 1 if the item can be reserved and 0 otherwise.
  // 
  function bit can_reserve(T item_to_reserve, bit external_lock = 0);
    I int_item;
    bit result;
    alloc_policy.in_use = this.in_use;
    if (alloc_policy.converter == null) begin
      `uvm_error("ITEM_ALLOCATOR", "alloc_policy.converter is null. can not be used.")
        return 0;
    end
    import_in_use(external_lock);
    int_item = alloc_policy.converter.serialize(item_to_reserve);
    result = alloc_policy.randomize(null) with {item == int_item;};
    done_in_use(external_lock);
    return result;
  endfunction: can_reserve

  // Function: reserve_item
  //
  // Reserve the specified ~item_to_reserve~.
  //
  // Return 1 if the item was successfully reserved
  // and 0 otherwise.
  function bit reserve_item(T item_to_reserve, bit external_lock = 0);
    I int_item;
    bit result;

    result = 0;
    alloc_policy.in_use = this.in_use;
    if (alloc_policy.converter == null) begin
      `uvm_error("ITEM_ALLOCATOR", "alloc_policy.converter is null. can not be used.")
      return 0;
    end
    import_in_use(external_lock);
    int_item = alloc_policy.converter.serialize(item_to_reserve);
    if (alloc_policy.randomize() with {item==int_item;})
      begin
        result = 1;

        this.in_use.push_back(alloc_policy.item);
        export_in_use(external_lock);
      end
    else
    begin
      done_in_use(external_lock);
      `uvm_error("ITEM-ALLOCATOR", $sformatf("Can not reserve item %d",item_to_reserve) )
    end
    return result;
  endfunction: reserve_item
  
  // Function: can_request
  //
  // Check if an item can be requsted according to specified ~alloc~ policy
  // Return 1 if the item can be requested and 0 otherwise.
  // 
  function bit can_request(input uvm_item_alloc_policy#(T, I) alloc = null, 
                           bit external_lock = 0);
    bit result;
    result = 0;
    
    if (alloc == null)
       alloc = alloc_policy;

    import_in_use(external_lock);
    alloc.in_use = this.in_use;
    result = alloc_policy.randomize(null);
    done_in_use(external_lock);
    return result;
  endfunction: can_request
  
  // Function: request_item
  //
  // Request and reserve an item accirding to specified ~alloc~ policy
  //
  // Return 1 if the item was successfully reserved
  // and to 0 otherwise.
  // output ~item~ is set to the allocated item, if allocation was successfull

  function bit request_item(uvm_item_alloc_policy#(T, I) alloc, 
                            output T item, input bit external_lock=0);
    bit result;
    result = 0;

    if (alloc == null)
      alloc = alloc_policy;

    import_in_use(external_lock);
    alloc.in_use = this.in_use;
    result = alloc.randomize();

    if (result) begin
      item = alloc.object;
      this.in_use.push_back(alloc.item);
      export_in_use(external_lock);
    end
    else begin
      done_in_use(external_lock);
      `uvm_error("ITEM-ALLOCATOR", "Can not request item" )
    end
    return result;
  endfunction: request_item
  
  // Function: release_item
  //
  // Release specified ~object~.
  //
  function void release_item(T object, bit external_lock = 0);
    I item;
    if (alloc_policy.converter == null) begin
      `uvm_error("ITEM_ALLOCATOR", "coverter is not set. can not be used")
      return;
    end
    item = alloc_policy.converter.serialize(object);
    import_in_use(external_lock);
    foreach (this.in_use[i]) begin
      if (this.in_use[i] == item) begin
        this.in_use.delete(i);
        export_in_use(external_lock);
        return;
      end
    end
    done_in_use(external_lock);
   `uvm_error("ITEM-ALLOCATOR", $sformatf("can not release item %0d. it is not currently allocated", item))
  endfunction: release_item
  
  // Function: release_all_items
  //
  // Release all currenly allocated items
  //
  function void release_all_items(bit external_lock = 0);
    start_in_use(external_lock);
    in_use.delete();
    export_in_use(external_lock);
  endfunction: release_all_items
  
  
   // Function: convert2string
   //
   // Create a human-readable description the currently allocated items.
   // 
  function string convert2string();
    string result;
    import_in_use(1); // do we need a task version of this function, which actually waits for lock?
    result = "Allocated items: \n";
    foreach (this.in_use[i]) begin
      $sformat(result, "%s   %0d", result,
               this.in_use[i]);
    end
    result = {result, "\n"};
    done_in_use(1);
    return result;
  endfunction: convert2string

endclass: uvm_item_allocator

`endif // ifndef UVM_ITEM_ALLOCATOR__SVH
