../08passive_ending/uvm_phase_objection.svh