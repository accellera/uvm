//----------------------------------------------------------------------
//   Copyright 2013 Freescale Semiconductor, Inc.
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------

program top;

import uvm_pkg::*;
`include "uvm_macros.svh"


class test extends uvm_test;

   `uvm_component_utils(test)

   function new(string name, uvm_component parent = null);
      super.new(name, parent);
   endfunction: new

   virtual task run();
      uvm_top.stop_request();
   endtask: run

   virtual function void report();
     int weight[20];
     int temp;
     uvm_dynamic_range_constraint#("RANDINT1") drc  = uvm_dynamic_range_constraint#("RANDINT1")::get_inst() ;
     uvm_dynamic_range_constraint#("RANDINT2") drc2 = uvm_dynamic_range_constraint#("RANDINT2")::get_inst() ;
     uvm_dynamic_range_constraint#("RANDINT3") drc3 = uvm_dynamic_range_constraint#("RANDINT3")::get_inst() ;
     uvm_dynamic_range_constraint#("RANDINT4") drc4 = uvm_dynamic_range_constraint#("RANDINT4")::get_inst() ;
     for(int unsigned index = 0; index != 100; ++index)
     begin
       temp = uvm_dynamic_range_constraint#("RANDINT1")::get_rand_value();
       weight[temp]++;
     end
     $write("Statistics for 100 randomizations of constraint RANDINT1:\n");
     for (int unsigned index=1; index != 20; ++index)
     begin
       $write("  %0d was chosen %0d times\n", index, weight[index]);
     end  
     
     $write("\n** UVM TEST PASSED **\n");
   endfunction: report

endclass: test

initial run_test();

endprogram: top
