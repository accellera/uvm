package mem_sequences;

  import uvm_pkg::*;
  import mem_agent::*;
  `include "uvm_macros.svh"

  `include "mem_sequences.svh"

endpackage