//----------------------------------------------------------------------
//   Copyright 2010 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------

//----------------------------------------------------------------------
// Generic Payload
//----------------------------------------------------------------------

`define ADDR_SIZE 64
const int unsigned addr_size = `ADDR_SIZE;
typedef bit[`ADDR_SIZE-1:0] tlm2_addr_t;

typedef enum
{
    TLM_READ_COMMAND,
    TLM_WRITE_COMMAND,
    TLM_IGNORE_COMMAND
} tlm_command_e;

typedef enum
{
    TLM_OK_RESPONSE = 1,
    TLM_INCOMPLETE_RESPONSE = 0,
    TLM_GENERIC_ERROR_RESPONSE = -1,
    TLM_ADDRESS_ERROR_RESPONSE = -2,
    TLM_COMMAND_ERROR_RESPONSE = -3,
    TLM_BURST_ERROR_RESPONSE = -4,
    TLM_BYTE_ENABLE_ERROR_RESPONSE = -5
} tlm_response_status_e;

//----------------------------------------------------------------------
// tlm2_generic_payload
//----------------------------------------------------------------------
virtual class tlm2_generic_payload extends uvm_sequence_item;

    local tlm2_addr_t            m_address;
    local tlm_command_e          m_command;
    local byte                   m_data[];
    local int unsigned           m_length;
    tlm_response_status_e  m_response_status;
    local bit                    m_dmi;
    local byte                   m_byte_enable[];
    local int unsigned           m_byte_enable_length;
    local int unsigned           m_streaming_width;

  function new(string name="");
    super.new(name);
    m_address = 0;
    m_command = TLM_IGNORE_COMMAND;
    m_length = 0;
    m_response_status = TLM_INCOMPLETE_RESPONSE;
    m_dmi = 0;
    m_byte_enable_length = 0;
    m_streaming_width = 0;
  endfunction

  function string convert2string();

    string msg;
    string addr_fmt;
    string s;
    int unsigned addr_chars = (addr_size >> 2) + ((addr_size & 'hf) > 0);

    $sformat(addr_fmt, "%%%0dx", addr_chars);
    $sformat(s, addr_fmt, m_address);
    $sformat(msg, "%s [%s] =", m_command.name(), s);

    for(int unsigned i = 0; i < m_data.size(); i++) begin
      $sformat(s, " %02x", m_data[i]);
      msg = { msg , s };
    end

    if(m_response_status != TLM_INCOMPLETE_RESPONSE)
      msg = { msg, " <-- ", get_response_string() };

    return msg;

  endfunction

  function void do_copy(uvm_object rhs);

    tlm2_generic_payload t;

    super.do_copy(rhs);

    if(rhs == null)
      return;
    if(!$cast(t, rhs))
      return;

    m_address            = t.m_address;
    m_command            = t.m_command;
    m_length             = t.m_length;
    m_response_status    = t.m_response_status;
    m_dmi                = t.m_dmi;
    m_byte_enable_length = t.m_byte_enable_length;
    m_streaming_width    = t.m_streaming_width;
    m_data               = t.m_data;
    m_byte_enable        = t.m_byte_enable;
  endfunction

  function uvm_object clone();
    tlm2_generic_payload t = new();
    t.copy(this);
    return t;
  endfunction

  // return an abbreviated response string
  function string get_response_string();

    case(m_response_status)
      TLM_OK_RESPONSE:                return "OK";
      TLM_INCOMPLETE_RESPONSE:        return "INCOMPLETE";
      TLM_GENERIC_ERROR_RESPONSE:     return "GENERIC_ERROR";
      TLM_ADDRESS_ERROR_RESPONSE:     return "ADDRESS_ERROR";
      TLM_COMMAND_ERROR_RESPONSE:     return "COMMAND_ERROR";
      TLM_BURST_ERROR_RESPONSE:       return "BURST_ERROR";
      TLM_BYTE_ENABLE_ERROR_RESPONSE: return "BYTE_ENABLE_ERROR";
    endcase

    // we should never get here
    return "UNKNOWN_RESPONSE";

  endfunction

  // accessors

  // command
  virtual function tlm_command_e get_command();
    return m_command;
  endfunction

  virtual function void set_command(tlm_command_e command);
    m_command = command;
  endfunction

  virtual function bit is_read();
    return (m_command == TLM_READ_COMMAND);
  endfunction

  virtual function void set_read();
    set_command(TLM_READ_COMMAND);
  endfunction

  virtual function bit is_write();
    return (m_command == TLM_WRITE_COMMAND);
  endfunction

  virtual function void set_write();
    set_command(TLM_WRITE_COMMAND);
  endfunction
  
  // address
  virtual function void set_address(tlm2_addr_t addr);
    m_address = addr;
  endfunction

  virtual function tlm2_addr_t get_address();
    return m_address;
  endfunction

  virtual function void get_data (output byte p []);
    p = m_data;
  endfunction

  virtual function void set_data_ptr(ref byte p []);
    m_data = p;
  endfunction

  virtual function int unsigned get_data_length();
    return m_length;
  endfunction

  virtual function void set_data_length(int unsigned length);
    m_length = length;
  endfunction

  virtual function int unsigned get_streaming_width();
    return m_streaming_width;
  endfunction

  virtual function void set_streaming_width(int unsigned width);
    m_streaming_width = width;
  endfunction

  virtual function void get_byte_enable(output byte p[]);
    p = m_byte_enable;
  endfunction

  virtual function void set_byte_enable(ref byte p[]);
    m_byte_enable = p;
  endfunction

  virtual function int unsigned get_byte_enable_length();
    return m_byte_enable_length;
  endfunction

  virtual function void set_byte_enable_length(int unsigned length);
    m_byte_enable_length = length;
  endfunction

 // DMI hint void set_dmi_allowed( bool );
  virtual function void set_dmi_allowed(bit dmi);
    m_dmi = dmi;
  endfunction

  virtual function bit is_dmi_allowed();
    return m_dmi;
  endfunction

// tlm_response_status get_response_status() const;
// void set_response_status( const tlm_response_status );
// std::string get_response_string();
// bool is_response_ok();
// bool is_response_error();

    
endclass

