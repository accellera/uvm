//----------------------------------------------------------------------
//   Copyright 2010 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------

//----------------------------------------------------------------------
// tlm2 package
//----------------------------------------------------------------------
package tlm2_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "tlm2_defines.svh"
  `include "tlm2_generic_payload.svh"
  `include "tlm2_ifs.svh"
  `include "tlm2_imps.svh"
  `include "tlm2_ports.svh"
  `include "tlm2_exports.svh"
  `include "tlm2_sockets_base.svh"
  `include "tlm2_sockets.svh"
  `include "tlm2_quantumkeeper.svh"
  `include "tlm2_peq.svh"

endpackage
