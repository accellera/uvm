package checker_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "checker.svh"

endpackage
