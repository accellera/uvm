//
//------------------------------------------------------------------------------
//   Copyright 2011 (Authors)
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------------------------

//Common testbench for these test case
//3.4        Advanced phase control 5
//  3.4.1         Killing phases. 5
//  3.4.2         Rerunning phases. 5
//  3.4.3         Fast-forwarding. 5

`include "top_uvc.svh"
`include "bot_uvc.svh"
`include "my_seqr.svh"

`include "test_base.svh"
