// $Id: methodology_noparm.svh,v 1.6 2009/05/12 21:02:29 redelman Exp $
//------------------------------------------------------------------------------
//   Copyright 2007-2009 Mentor Graphics Corporation
//   Copyright 2007-2009 Cadence Design Systems, Inc.
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------------------------

`ifndef UVM_METH_SVH
`define UVM_METH_SVH

  `include "methodology/sequences/uvm_sequence_item.svh"
  `include "methodology/sequences/uvm_sequencer_base.svh"
  `include "methodology/sequences/uvm_sequence_base.svh"

  `include "methodology/uvm_meth_defines.svh"

  `include "methodology/uvm_monitor.svh"
  `include "methodology/uvm_scoreboard.svh" 
  `include "methodology/uvm_agent.svh"
  `include "methodology/uvm_env.svh"
  `include "methodology/uvm_test.svh"

`endif //UVM_METH_SVH
