// test

