program top;

import uvm_pkg::*;
`include "uvm_macros.svh"

class test extends uvm_test;

   `uvm_component_utils(test)

   function new(string name, uvm_component parent);
      super.new(name, parent);
   endfunction

   task run();
     for (int i = 0; i < 20; i++) begin
       #100;
       `uvm_error("TESTERR", "An error.")
     end
   endtask

endclass


initial
  begin
     run_test();
  end

final
  begin
    if ($time == 300)
      $write("UVM TEST EXPECT 3 UVM_ERROR\n");
      $write("** UVM TEST PASSED **\n");
  end

endprogram
